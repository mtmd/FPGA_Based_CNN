`ifndef _parameters_vh
`define _parameters_vh
`define START				1
`define CHECK_OUTPUT		2
`define CHECK_OFM			3
`define CHECK_IFM			4
`define CHECK_WEIGHT		5
`define CHECK_RESULT		6
`define CHECK_LOOPS		8
`define CHECK_WB			7
`endif