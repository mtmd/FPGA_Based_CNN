module clock (
input clk_in,
output clk_out

);
assign clk_out = clk_in;
endmodule